// Benchmark "AddressGenerator_4096_pe1" written by ABC on Sat Mar 13 15:56:33 2021

module AddressGenerator_4096_pe1 ( 
    inp13, inp12, inp11, inp10, inp9, inp8, inp7, inp6, inp5, inp4, inp3,
    inp2, inp1, inp0,
    otp43, otp42, otp41, otp40, otp39, otp38, otp37, otp36, otp35, otp34,
    otp33, otp32, otp31, otp30, otp29, otp28, otp27, otp26, otp25, otp24,
    otp23, otp22, otp21, otp20, otp19, otp18, otp17, otp16, otp15, otp14,
    otp13, otp12, otp11, otp10, otp9, otp8, otp7, otp6, otp5, otp4, otp3,
    otp2, otp1, otp0  );
  input  inp13, inp12, inp11, inp10, inp9, inp8, inp7, inp6, inp5, inp4,
    inp3, inp2, inp1, inp0;
  output otp43, otp42, otp41, otp40, otp39, otp38, otp37, otp36, otp35, otp34,
    otp33, otp32, otp31, otp30, otp29, otp28, otp27, otp26, otp25, otp24,
    otp23, otp22, otp21, otp20, otp19, otp18, otp17, otp16, otp15, otp14,
    otp13, otp12, otp11, otp10, otp9, otp8, otp7, otp6, otp5, otp4, otp3,
    otp2, otp1, otp0;
  wire new_n59_, new_n60_, new_n61_, new_n62_, new_n63_, new_n64_, new_n65_,
    new_n66_, new_n67_, new_n68_, new_n69_, new_n70_, new_n71_, new_n72_,
    new_n73_, new_n74_, new_n75_, new_n76_, new_n77_, new_n78_, new_n79_,
    new_n80_, new_n81_, new_n82_, new_n83_, new_n84_, new_n85_, new_n86_,
    new_n87_, new_n88_, new_n89_, new_n90_, new_n91_, new_n92_, new_n93_,
    new_n94_, new_n95_, new_n96_, new_n97_, new_n98_, new_n99_, new_n100_,
    new_n101_, new_n102_, new_n103_, new_n104_, new_n105_, new_n106_,
    new_n107_, new_n108_, new_n109_, new_n110_, new_n111_, new_n112_,
    new_n113_, new_n114_, new_n115_, new_n116_, new_n117_, new_n118_,
    new_n119_, new_n120_, new_n121_, new_n122_, new_n123_, new_n124_,
    new_n125_, new_n126_, new_n127_, new_n128_, new_n129_, new_n130_,
    new_n131_, new_n132_, new_n133_, new_n134_, new_n135_, new_n136_,
    new_n137_, new_n138_, new_n139_, new_n140_, new_n141_, new_n142_,
    new_n143_, new_n144_, new_n145_, new_n146_, new_n147_, new_n148_,
    new_n149_, new_n150_, new_n151_, new_n152_, new_n154_, new_n155_,
    new_n156_, new_n157_, new_n158_, new_n159_, new_n160_, new_n161_,
    new_n163_, new_n164_, new_n165_, new_n166_, new_n167_, new_n168_,
    new_n169_, new_n170_, new_n171_, new_n172_, new_n173_, new_n174_,
    new_n175_, new_n176_, new_n177_, new_n178_, new_n179_, new_n180_,
    new_n181_, new_n182_, new_n183_, new_n184_, new_n185_, new_n186_,
    new_n187_, new_n188_, new_n189_, new_n190_, new_n191_, new_n192_,
    new_n193_, new_n194_, new_n195_, new_n196_, new_n197_, new_n198_,
    new_n199_, new_n200_, new_n201_, new_n202_, new_n203_, new_n204_,
    new_n205_, new_n206_, new_n207_, new_n208_, new_n209_, new_n210_,
    new_n211_, new_n212_, new_n213_, new_n214_, new_n215_, new_n216_,
    new_n217_, new_n218_, new_n219_, new_n220_, new_n221_, new_n222_,
    new_n223_, new_n224_, new_n225_, new_n226_, new_n227_, new_n228_,
    new_n229_, new_n230_, new_n231_, new_n232_, new_n233_, new_n234_,
    new_n235_, new_n236_, new_n237_, new_n238_, new_n239_, new_n240_,
    new_n241_, new_n242_, new_n243_, new_n244_, new_n245_, new_n246_,
    new_n248_, new_n249_, new_n250_, new_n251_, new_n252_, new_n253_,
    new_n254_, new_n255_, new_n256_, new_n257_, new_n258_, new_n259_,
    new_n260_, new_n261_, new_n262_, new_n263_, new_n264_, new_n265_,
    new_n266_, new_n267_, new_n268_, new_n269_, new_n270_, new_n271_,
    new_n272_, new_n273_, new_n274_, new_n275_, new_n276_, new_n277_,
    new_n278_, new_n279_, new_n280_, new_n281_, new_n282_, new_n283_,
    new_n284_, new_n285_, new_n286_, new_n287_, new_n288_, new_n289_,
    new_n290_, new_n291_, new_n292_, new_n293_, new_n294_, new_n295_,
    new_n296_, new_n297_, new_n298_, new_n299_, new_n300_, new_n301_,
    new_n302_, new_n304_, new_n305_, new_n306_, new_n307_, new_n308_,
    new_n309_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n317_, new_n318_, new_n319_, new_n320_, new_n321_, new_n322_,
    new_n323_, new_n325_, new_n326_, new_n327_, new_n329_, new_n330_,
    new_n331_, new_n332_, new_n333_, new_n334_, new_n335_, new_n336_,
    new_n337_, new_n338_, new_n339_, new_n341_, new_n342_, new_n343_,
    new_n344_, new_n345_, new_n346_, new_n347_, new_n348_, new_n350_,
    new_n351_, new_n352_, new_n353_, new_n354_, new_n355_, new_n356_,
    new_n357_, new_n358_, new_n359_, new_n360_, new_n361_, new_n362_,
    new_n363_, new_n364_, new_n365_, new_n366_, new_n367_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n375_, new_n376_,
    new_n377_, new_n378_, new_n379_, new_n380_, new_n381_, new_n382_,
    new_n383_, new_n384_, new_n385_, new_n386_, new_n387_, new_n388_,
    new_n389_, new_n390_, new_n391_, new_n392_, new_n393_, new_n394_,
    new_n396_, new_n397_, new_n398_, new_n399_, new_n400_, new_n401_,
    new_n402_, new_n405_, new_n407_, new_n409_, new_n411_, new_n412_,
    new_n413_, new_n415_, new_n417_, new_n418_, new_n419_, new_n421_,
    new_n423_, new_n424_, new_n425_, new_n426_, new_n427_, new_n429_,
    new_n431_, new_n432_, new_n433_, new_n434_, new_n435_, new_n436_,
    new_n437_, new_n438_, new_n439_, new_n441_, new_n442_, new_n443_,
    new_n444_, new_n445_, new_n446_, new_n447_, new_n448_, new_n449_,
    new_n450_, new_n451_, new_n452_, new_n453_, new_n454_, new_n455_,
    new_n457_, new_n458_, new_n459_, new_n460_, new_n461_, new_n462_,
    new_n463_, new_n464_, new_n465_, new_n466_, new_n467_, new_n468_,
    new_n469_, new_n470_, new_n471_, new_n472_, new_n473_, new_n474_,
    new_n475_, new_n476_, new_n477_, new_n478_, new_n479_, new_n481_,
    new_n482_, new_n483_, new_n484_, new_n485_, new_n486_, new_n487_,
    new_n488_, new_n489_, new_n490_, new_n491_, new_n492_, new_n494_,
    new_n495_, new_n496_, new_n497_, new_n498_, new_n499_, new_n500_,
    new_n501_, new_n502_, new_n503_, new_n504_, new_n505_, new_n506_,
    new_n507_, new_n508_, new_n509_, new_n510_, new_n511_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n523_, new_n524_, new_n525_, new_n526_,
    new_n527_, new_n528_, new_n529_, new_n530_, new_n531_, new_n532_,
    new_n533_, new_n534_, new_n536_, new_n537_, new_n538_, new_n539_,
    new_n540_, new_n541_, new_n542_, new_n543_, new_n544_, new_n545_,
    new_n546_, new_n547_, new_n548_, new_n549_, new_n550_, new_n551_,
    new_n553_, new_n554_, new_n555_, new_n556_, new_n557_, new_n558_,
    new_n559_, new_n560_, new_n561_, new_n562_, new_n563_, new_n564_,
    new_n565_, new_n566_, new_n567_, new_n568_, new_n569_, new_n570_,
    new_n571_, new_n572_, new_n573_, new_n574_, new_n576_, new_n578_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n593_,
    new_n595_, new_n596_, new_n597_, new_n598_, new_n599_, new_n600_,
    new_n601_, new_n602_, new_n603_, new_n604_, new_n605_, new_n606_,
    new_n608_, new_n609_, new_n610_, new_n612_, new_n613_, new_n614_,
    new_n615_, new_n616_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_;
  assign new_n59_ = ~inp13 & ~inp12;
  assign new_n60_ = inp9 & inp8;
  assign new_n61_ = ~inp9 & ~inp8;
  assign new_n62_ = ~new_n60_ & ~new_n61_;
  assign new_n63_ = inp11 & ~inp10;
  assign new_n64_ = inp7 & new_n63_;
  assign new_n65_ = inp11 & inp10;
  assign new_n66_ = inp7 & ~inp6;
  assign new_n67_ = ~inp7 & inp6;
  assign new_n68_ = ~new_n66_ & ~new_n67_;
  assign new_n69_ = new_n65_ & ~new_n68_;
  assign new_n70_ = ~new_n64_ & ~new_n69_;
  assign new_n71_ = ~inp11 & ~inp10;
  assign new_n72_ = new_n70_ & ~new_n71_;
  assign new_n73_ = ~new_n62_ & new_n72_;
  assign new_n74_ = new_n62_ & ~new_n70_;
  assign new_n75_ = ~inp9 & new_n71_;
  assign new_n76_ = ~new_n74_ & ~new_n75_;
  assign new_n77_ = ~new_n73_ & new_n76_;
  assign new_n78_ = new_n59_ & ~new_n77_;
  assign new_n79_ = inp9 & ~inp4;
  assign new_n80_ = ~inp9 & inp4;
  assign new_n81_ = ~new_n79_ & ~new_n80_;
  assign new_n82_ = inp2 & ~inp1;
  assign new_n83_ = ~inp2 & inp1;
  assign new_n84_ = ~new_n82_ & ~new_n83_;
  assign new_n85_ = inp0 & ~new_n84_;
  assign new_n86_ = ~inp0 & new_n84_;
  assign new_n87_ = ~new_n85_ & ~new_n86_;
  assign new_n88_ = ~inp3 & ~new_n87_;
  assign new_n89_ = inp3 & new_n87_;
  assign new_n90_ = ~new_n88_ & ~new_n89_;
  assign new_n91_ = ~new_n71_ & ~new_n90_;
  assign new_n92_ = inp3 & ~new_n84_;
  assign new_n93_ = ~inp3 & new_n84_;
  assign new_n94_ = ~new_n92_ & ~new_n93_;
  assign new_n95_ = ~inp11 & ~new_n94_;
  assign new_n96_ = ~inp10 & new_n95_;
  assign new_n97_ = ~new_n91_ & ~new_n96_;
  assign new_n98_ = ~inp12 & ~new_n97_;
  assign new_n99_ = inp13 & new_n98_;
  assign new_n100_ = inp10 & ~inp2;
  assign new_n101_ = ~new_n63_ & ~new_n100_;
  assign new_n102_ = ~inp3 & ~new_n101_;
  assign new_n103_ = inp3 & inp2;
  assign new_n104_ = inp11 & ~new_n103_;
  assign new_n105_ = inp10 & ~new_n104_;
  assign new_n106_ = ~new_n102_ & ~new_n105_;
  assign new_n107_ = inp12 & ~new_n106_;
  assign new_n108_ = ~inp13 & new_n107_;
  assign new_n109_ = ~new_n99_ & ~new_n108_;
  assign new_n110_ = ~new_n81_ & ~new_n109_;
  assign new_n111_ = ~inp13 & inp12;
  assign new_n112_ = inp9 & new_n71_;
  assign new_n113_ = new_n111_ & new_n112_;
  assign new_n114_ = ~inp3 & ~inp2;
  assign new_n115_ = ~new_n103_ & ~new_n114_;
  assign new_n116_ = new_n65_ & new_n111_;
  assign new_n117_ = new_n115_ & new_n116_;
  assign new_n118_ = new_n63_ & new_n111_;
  assign new_n119_ = inp3 & new_n118_;
  assign new_n120_ = ~new_n117_ & ~new_n119_;
  assign new_n121_ = inp1 & new_n71_;
  assign new_n122_ = ~inp1 & ~inp0;
  assign new_n123_ = inp1 & inp0;
  assign new_n124_ = ~new_n122_ & ~new_n123_;
  assign new_n125_ = ~new_n71_ & new_n124_;
  assign new_n126_ = ~new_n121_ & ~new_n125_;
  assign new_n127_ = new_n115_ & ~new_n126_;
  assign new_n128_ = inp13 & ~inp12;
  assign new_n129_ = ~new_n115_ & new_n126_;
  assign new_n130_ = new_n128_ & ~new_n129_;
  assign new_n131_ = ~new_n127_ & new_n130_;
  assign new_n132_ = new_n120_ & ~new_n131_;
  assign new_n133_ = new_n81_ & ~new_n132_;
  assign new_n134_ = ~new_n113_ & ~new_n133_;
  assign new_n135_ = ~new_n110_ & new_n134_;
  assign new_n136_ = inp6 & ~inp5;
  assign new_n137_ = ~inp6 & inp5;
  assign new_n138_ = ~new_n136_ & ~new_n137_;
  assign new_n139_ = ~inp8 & ~inp7;
  assign new_n140_ = inp8 & inp7;
  assign new_n141_ = ~new_n139_ & ~new_n140_;
  assign new_n142_ = new_n138_ & ~new_n141_;
  assign new_n143_ = ~new_n138_ & new_n141_;
  assign new_n144_ = ~new_n142_ & ~new_n143_;
  assign new_n145_ = ~new_n135_ & new_n144_;
  assign new_n146_ = new_n81_ & ~new_n109_;
  assign new_n147_ = new_n75_ & new_n111_;
  assign new_n148_ = ~new_n81_ & ~new_n132_;
  assign new_n149_ = ~new_n147_ & ~new_n148_;
  assign new_n150_ = ~new_n146_ & new_n149_;
  assign new_n151_ = ~new_n144_ & ~new_n150_;
  assign new_n152_ = ~new_n145_ & ~new_n151_;
  assign otp43 = new_n78_ | ~new_n152_;
  assign new_n154_ = new_n62_ & new_n72_;
  assign new_n155_ = ~new_n62_ & ~new_n70_;
  assign new_n156_ = ~new_n112_ & ~new_n155_;
  assign new_n157_ = ~new_n154_ & new_n156_;
  assign new_n158_ = new_n59_ & ~new_n157_;
  assign new_n159_ = new_n144_ & ~new_n150_;
  assign new_n160_ = ~new_n135_ & ~new_n144_;
  assign new_n161_ = ~new_n159_ & ~new_n160_;
  assign otp42 = new_n158_ | ~new_n161_;
  assign new_n163_ = inp10 & inp9;
  assign new_n164_ = ~inp13 & new_n163_;
  assign new_n165_ = ~inp12 & ~inp11;
  assign new_n166_ = ~new_n164_ & new_n165_;
  assign new_n167_ = inp10 & inp1;
  assign new_n168_ = ~inp5 & ~inp4;
  assign new_n169_ = inp5 & inp4;
  assign new_n170_ = ~new_n168_ & ~new_n169_;
  assign new_n171_ = new_n115_ & ~new_n170_;
  assign new_n172_ = ~new_n115_ & new_n170_;
  assign new_n173_ = ~new_n171_ & ~new_n172_;
  assign new_n174_ = ~new_n167_ & ~new_n173_;
  assign new_n175_ = new_n167_ & new_n173_;
  assign new_n176_ = ~new_n174_ & ~new_n175_;
  assign new_n177_ = ~new_n62_ & new_n68_;
  assign new_n178_ = new_n62_ & ~new_n68_;
  assign new_n179_ = ~new_n177_ & ~new_n178_;
  assign new_n180_ = ~new_n176_ & new_n179_;
  assign new_n181_ = new_n176_ & ~new_n179_;
  assign new_n182_ = inp13 & ~new_n181_;
  assign new_n183_ = ~new_n180_ & new_n182_;
  assign new_n184_ = new_n166_ & ~new_n183_;
  assign new_n185_ = new_n115_ & ~new_n124_;
  assign new_n186_ = ~new_n115_ & new_n124_;
  assign new_n187_ = ~new_n185_ & ~new_n186_;
  assign new_n188_ = new_n128_ & ~new_n187_;
  assign new_n189_ = inp10 & inp3;
  assign new_n190_ = new_n111_ & new_n189_;
  assign new_n191_ = ~new_n188_ & ~new_n190_;
  assign new_n192_ = new_n179_ & ~new_n191_;
  assign new_n193_ = ~new_n170_ & new_n192_;
  assign new_n194_ = new_n111_ & ~new_n189_;
  assign new_n195_ = new_n128_ & new_n187_;
  assign new_n196_ = ~new_n194_ & ~new_n195_;
  assign new_n197_ = new_n170_ & new_n179_;
  assign new_n198_ = ~new_n196_ & new_n197_;
  assign new_n199_ = new_n170_ & new_n191_;
  assign new_n200_ = ~new_n170_ & new_n196_;
  assign new_n201_ = ~new_n199_ & ~new_n200_;
  assign new_n202_ = ~new_n179_ & new_n201_;
  assign new_n203_ = inp10 & inp7;
  assign new_n204_ = ~new_n62_ & ~new_n203_;
  assign new_n205_ = new_n62_ & new_n203_;
  assign new_n206_ = ~new_n204_ & ~new_n205_;
  assign new_n207_ = new_n59_ & ~new_n206_;
  assign new_n208_ = ~new_n202_ & ~new_n207_;
  assign new_n209_ = ~new_n198_ & new_n208_;
  assign new_n210_ = ~new_n193_ & new_n209_;
  assign new_n211_ = inp11 & ~new_n210_;
  assign new_n212_ = inp8 & ~inp5;
  assign new_n213_ = ~inp8 & inp5;
  assign new_n214_ = ~new_n212_ & ~new_n213_;
  assign new_n215_ = ~inp10 & ~inp4;
  assign new_n216_ = inp10 & inp4;
  assign new_n217_ = ~new_n215_ & ~new_n216_;
  assign new_n218_ = ~new_n187_ & new_n217_;
  assign new_n219_ = new_n187_ & ~new_n217_;
  assign new_n220_ = inp13 & ~new_n219_;
  assign new_n221_ = ~new_n218_ & new_n220_;
  assign new_n222_ = ~inp13 & ~inp10;
  assign new_n223_ = ~new_n221_ & ~new_n222_;
  assign new_n224_ = ~new_n214_ & new_n223_;
  assign new_n225_ = ~inp9 & new_n224_;
  assign new_n226_ = ~inp9 & new_n221_;
  assign new_n227_ = ~new_n164_ & ~new_n226_;
  assign new_n228_ = new_n214_ & ~new_n227_;
  assign new_n229_ = new_n62_ & new_n222_;
  assign new_n230_ = ~new_n228_ & ~new_n229_;
  assign new_n231_ = ~new_n225_ & new_n230_;
  assign new_n232_ = ~new_n68_ & new_n231_;
  assign new_n233_ = inp12 & ~inp11;
  assign new_n234_ = new_n214_ & new_n223_;
  assign new_n235_ = ~inp8 & new_n222_;
  assign new_n236_ = ~inp9 & ~new_n235_;
  assign new_n237_ = ~new_n234_ & new_n236_;
  assign new_n238_ = inp8 & new_n222_;
  assign new_n239_ = inp9 & ~new_n238_;
  assign new_n240_ = ~new_n237_ & ~new_n239_;
  assign new_n241_ = ~new_n214_ & ~new_n227_;
  assign new_n242_ = new_n68_ & ~new_n241_;
  assign new_n243_ = ~new_n240_ & new_n242_;
  assign new_n244_ = new_n233_ & ~new_n243_;
  assign new_n245_ = ~new_n232_ & new_n244_;
  assign new_n246_ = ~new_n211_ & ~new_n245_;
  assign otp41 = new_n184_ | ~new_n246_;
  assign new_n248_ = inp11 & ~new_n196_;
  assign new_n249_ = new_n115_ & ~new_n167_;
  assign new_n250_ = ~new_n115_ & new_n167_;
  assign new_n251_ = ~new_n249_ & ~new_n250_;
  assign new_n252_ = new_n128_ & new_n251_;
  assign new_n253_ = ~inp11 & new_n252_;
  assign new_n254_ = new_n170_ & ~new_n253_;
  assign new_n255_ = ~new_n248_ & new_n254_;
  assign new_n256_ = inp11 & new_n190_;
  assign new_n257_ = ~inp11 & new_n167_;
  assign new_n258_ = inp11 & new_n124_;
  assign new_n259_ = ~new_n257_ & ~new_n258_;
  assign new_n260_ = ~new_n115_ & new_n259_;
  assign new_n261_ = new_n115_ & ~new_n259_;
  assign new_n262_ = new_n128_ & ~new_n261_;
  assign new_n263_ = ~new_n260_ & new_n262_;
  assign new_n264_ = ~new_n256_ & ~new_n263_;
  assign new_n265_ = ~new_n170_ & new_n264_;
  assign new_n266_ = ~new_n255_ & ~new_n265_;
  assign new_n267_ = inp10 & inp5;
  assign new_n268_ = ~inp11 & new_n267_;
  assign new_n269_ = new_n111_ & new_n268_;
  assign new_n270_ = ~new_n266_ & ~new_n269_;
  assign new_n271_ = ~new_n179_ & ~new_n270_;
  assign new_n272_ = inp13 & inp12;
  assign new_n273_ = ~inp9 & new_n272_;
  assign new_n274_ = ~new_n170_ & new_n187_;
  assign new_n275_ = new_n170_ & ~new_n187_;
  assign new_n276_ = ~new_n274_ & ~new_n275_;
  assign new_n277_ = ~inp10 & ~inp8;
  assign new_n278_ = inp10 & inp8;
  assign new_n279_ = ~new_n277_ & ~new_n278_;
  assign new_n280_ = new_n68_ & ~new_n279_;
  assign new_n281_ = ~new_n68_ & new_n279_;
  assign new_n282_ = ~new_n280_ & ~new_n281_;
  assign new_n283_ = ~new_n276_ & ~new_n282_;
  assign new_n284_ = new_n276_ & new_n282_;
  assign new_n285_ = ~new_n283_ & ~new_n284_;
  assign new_n286_ = new_n273_ & new_n285_;
  assign new_n287_ = new_n59_ & new_n163_;
  assign new_n288_ = ~new_n286_ & ~new_n287_;
  assign new_n289_ = new_n111_ & ~new_n267_;
  assign new_n290_ = new_n128_ & new_n176_;
  assign new_n291_ = ~new_n289_ & ~new_n290_;
  assign new_n292_ = new_n179_ & ~new_n291_;
  assign new_n293_ = ~inp11 & ~new_n292_;
  assign new_n294_ = new_n288_ & new_n293_;
  assign new_n295_ = new_n179_ & new_n201_;
  assign new_n296_ = inp11 & ~new_n295_;
  assign new_n297_ = new_n62_ & ~new_n203_;
  assign new_n298_ = ~new_n62_ & new_n203_;
  assign new_n299_ = ~new_n297_ & ~new_n298_;
  assign new_n300_ = new_n59_ & ~new_n299_;
  assign new_n301_ = new_n296_ & ~new_n300_;
  assign new_n302_ = ~new_n294_ & ~new_n301_;
  assign otp40 = new_n271_ | new_n302_;
  assign new_n304_ = ~inp10 & new_n165_;
  assign new_n305_ = ~inp9 & ~new_n304_;
  assign new_n306_ = ~inp12 & new_n112_;
  assign new_n307_ = ~new_n305_ & ~new_n306_;
  assign new_n308_ = ~inp13 & ~new_n307_;
  assign new_n309_ = ~inp9 & new_n128_;
  assign otp39 = new_n308_ | new_n309_;
  assign new_n311_ = ~inp11 & new_n59_;
  assign new_n312_ = ~new_n272_ & ~new_n311_;
  assign new_n313_ = ~new_n62_ & new_n312_;
  assign new_n314_ = inp8 & new_n59_;
  assign new_n315_ = ~inp11 & new_n314_;
  assign otp38 = new_n313_ | new_n315_;
  assign new_n317_ = new_n59_ & ~new_n65_;
  assign new_n318_ = ~new_n272_ & ~new_n317_;
  assign new_n319_ = ~inp9 & ~new_n141_;
  assign new_n320_ = inp9 & new_n141_;
  assign new_n321_ = ~new_n319_ & ~new_n320_;
  assign new_n322_ = new_n318_ & ~new_n321_;
  assign new_n323_ = inp7 & new_n317_;
  assign otp37 = new_n322_ | new_n323_;
  assign new_n325_ = inp6 & new_n59_;
  assign new_n326_ = ~new_n111_ & ~new_n128_;
  assign new_n327_ = ~new_n179_ & ~new_n326_;
  assign otp36 = new_n325_ | new_n327_;
  assign new_n329_ = inp12 & ~new_n71_;
  assign new_n330_ = inp5 & ~new_n329_;
  assign new_n331_ = ~inp13 & new_n330_;
  assign new_n332_ = ~inp13 & ~new_n71_;
  assign new_n333_ = inp12 & ~new_n332_;
  assign new_n334_ = ~new_n59_ & ~new_n333_;
  assign new_n335_ = ~new_n321_ & new_n334_;
  assign new_n336_ = new_n138_ & new_n335_;
  assign new_n337_ = new_n321_ & new_n334_;
  assign new_n338_ = ~new_n138_ & new_n337_;
  assign new_n339_ = ~new_n336_ & ~new_n338_;
  assign otp35 = new_n331_ | ~new_n339_;
  assign new_n341_ = inp12 & inp11;
  assign new_n342_ = ~inp13 & inp4;
  assign new_n343_ = ~new_n341_ & new_n342_;
  assign new_n344_ = ~inp13 & new_n341_;
  assign new_n345_ = ~new_n128_ & ~new_n344_;
  assign new_n346_ = ~new_n170_ & ~new_n179_;
  assign new_n347_ = ~new_n197_ & ~new_n346_;
  assign new_n348_ = ~new_n345_ & ~new_n347_;
  assign otp34 = new_n343_ | new_n348_;
  assign new_n350_ = inp4 & ~inp3;
  assign new_n351_ = ~inp4 & inp3;
  assign new_n352_ = ~new_n350_ & ~new_n351_;
  assign new_n353_ = ~new_n116_ & ~new_n128_;
  assign new_n354_ = new_n321_ & ~new_n353_;
  assign new_n355_ = ~new_n138_ & ~new_n354_;
  assign new_n356_ = ~new_n321_ & ~new_n353_;
  assign new_n357_ = new_n138_ & ~new_n356_;
  assign new_n358_ = ~new_n355_ & ~new_n357_;
  assign new_n359_ = new_n352_ & new_n358_;
  assign new_n360_ = inp12 & new_n65_;
  assign new_n361_ = ~inp13 & inp3;
  assign new_n362_ = ~new_n360_ & new_n361_;
  assign new_n363_ = ~new_n138_ & ~new_n356_;
  assign new_n364_ = new_n138_ & ~new_n354_;
  assign new_n365_ = ~new_n363_ & ~new_n364_;
  assign new_n366_ = ~new_n352_ & new_n365_;
  assign new_n367_ = ~new_n362_ & ~new_n366_;
  assign otp33 = new_n359_ | ~new_n367_;
  assign new_n369_ = new_n173_ & ~new_n179_;
  assign new_n370_ = ~new_n173_ & new_n179_;
  assign new_n371_ = ~new_n369_ & ~new_n370_;
  assign new_n372_ = new_n128_ & ~new_n371_;
  assign new_n373_ = ~inp13 & inp2;
  assign otp32 = new_n372_ | new_n373_;
  assign new_n375_ = ~inp13 & inp1;
  assign new_n376_ = ~new_n71_ & ~new_n321_;
  assign new_n377_ = ~new_n138_ & ~new_n376_;
  assign new_n378_ = ~new_n71_ & new_n321_;
  assign new_n379_ = new_n138_ & ~new_n378_;
  assign new_n380_ = ~new_n377_ & ~new_n379_;
  assign new_n381_ = ~new_n352_ & ~new_n380_;
  assign new_n382_ = new_n138_ & ~new_n376_;
  assign new_n383_ = ~new_n138_ & ~new_n378_;
  assign new_n384_ = ~new_n382_ & ~new_n383_;
  assign new_n385_ = new_n352_ & ~new_n384_;
  assign new_n386_ = ~new_n381_ & ~new_n385_;
  assign new_n387_ = new_n84_ & new_n386_;
  assign new_n388_ = ~new_n352_ & ~new_n384_;
  assign new_n389_ = new_n352_ & ~new_n380_;
  assign new_n390_ = ~new_n388_ & ~new_n389_;
  assign new_n391_ = ~new_n84_ & new_n390_;
  assign new_n392_ = ~new_n121_ & ~new_n391_;
  assign new_n393_ = ~new_n387_ & new_n392_;
  assign new_n394_ = new_n128_ & ~new_n393_;
  assign otp31 = new_n375_ | new_n394_;
  assign new_n396_ = ~new_n179_ & new_n276_;
  assign new_n397_ = new_n179_ & ~new_n276_;
  assign new_n398_ = ~new_n396_ & ~new_n397_;
  assign new_n399_ = inp11 & new_n128_;
  assign new_n400_ = new_n398_ & new_n399_;
  assign new_n401_ = inp13 & ~new_n165_;
  assign new_n402_ = inp0 & ~new_n401_;
  assign otp30 = new_n400_ | new_n402_;
  assign otp29 = inp9 & ~new_n272_;
  assign new_n405_ = new_n62_ & new_n312_;
  assign otp28 = new_n315_ | new_n405_;
  assign new_n407_ = new_n318_ & new_n321_;
  assign otp27 = new_n323_ | new_n407_;
  assign new_n409_ = new_n179_ & ~new_n326_;
  assign otp26 = new_n325_ | new_n409_;
  assign new_n411_ = ~new_n138_ & new_n335_;
  assign new_n412_ = new_n138_ & new_n337_;
  assign new_n413_ = ~new_n411_ & ~new_n412_;
  assign otp25 = new_n331_ | ~new_n413_;
  assign new_n415_ = ~new_n345_ & new_n347_;
  assign otp24 = new_n343_ | new_n415_;
  assign new_n417_ = new_n352_ & new_n365_;
  assign new_n418_ = ~new_n352_ & new_n358_;
  assign new_n419_ = ~new_n362_ & ~new_n418_;
  assign otp23 = new_n417_ | ~new_n419_;
  assign new_n421_ = new_n128_ & new_n371_;
  assign otp22 = new_n373_ | new_n421_;
  assign new_n423_ = ~new_n84_ & new_n386_;
  assign new_n424_ = new_n84_ & new_n390_;
  assign new_n425_ = ~new_n121_ & ~new_n424_;
  assign new_n426_ = ~new_n423_ & new_n425_;
  assign new_n427_ = new_n128_ & ~new_n426_;
  assign otp21 = new_n375_ | new_n427_;
  assign new_n429_ = ~new_n398_ & new_n399_;
  assign otp20 = new_n402_ | new_n429_;
  assign new_n431_ = new_n59_ & ~new_n63_;
  assign new_n432_ = new_n233_ & new_n285_;
  assign new_n433_ = inp13 & ~new_n432_;
  assign new_n434_ = ~new_n431_ & ~new_n433_;
  assign new_n435_ = ~inp9 & new_n434_;
  assign new_n436_ = ~inp13 & new_n306_;
  assign new_n437_ = ~inp12 & ~inp9;
  assign new_n438_ = ~new_n222_ & new_n437_;
  assign new_n439_ = ~new_n436_ & ~new_n438_;
  assign otp19 = new_n435_ | ~new_n439_;
  assign new_n441_ = ~inp9 & new_n233_;
  assign new_n442_ = inp13 & new_n441_;
  assign new_n443_ = ~inp7 & ~new_n279_;
  assign new_n444_ = inp7 & new_n279_;
  assign new_n445_ = ~new_n443_ & ~new_n444_;
  assign new_n446_ = new_n84_ & new_n138_;
  assign new_n447_ = ~new_n84_ & ~new_n138_;
  assign new_n448_ = ~new_n446_ & ~new_n447_;
  assign new_n449_ = new_n352_ & ~new_n448_;
  assign new_n450_ = ~new_n352_ & new_n448_;
  assign new_n451_ = ~new_n449_ & ~new_n450_;
  assign new_n452_ = new_n445_ & ~new_n451_;
  assign new_n453_ = ~new_n445_ & new_n451_;
  assign new_n454_ = ~new_n452_ & ~new_n453_;
  assign new_n455_ = new_n442_ & ~new_n454_;
  assign otp18 = otp38 | new_n455_;
  assign new_n457_ = new_n65_ & ~new_n321_;
  assign new_n458_ = ~inp13 & ~new_n457_;
  assign new_n459_ = inp12 & new_n321_;
  assign new_n460_ = ~inp12 & ~inp7;
  assign new_n461_ = ~new_n65_ & ~new_n460_;
  assign new_n462_ = ~new_n459_ & new_n461_;
  assign new_n463_ = new_n458_ & ~new_n462_;
  assign new_n464_ = inp10 & ~inp6;
  assign new_n465_ = ~inp10 & inp6;
  assign new_n466_ = ~new_n464_ & ~new_n465_;
  assign new_n467_ = ~new_n173_ & new_n466_;
  assign new_n468_ = new_n173_ & ~new_n466_;
  assign new_n469_ = ~new_n467_ & ~new_n468_;
  assign new_n470_ = inp12 & new_n469_;
  assign new_n471_ = ~new_n341_ & ~new_n470_;
  assign new_n472_ = new_n319_ & new_n471_;
  assign new_n473_ = ~inp12 & new_n320_;
  assign new_n474_ = ~inp9 & new_n141_;
  assign new_n475_ = new_n233_ & new_n474_;
  assign new_n476_ = new_n469_ & new_n475_;
  assign new_n477_ = ~new_n473_ & ~new_n476_;
  assign new_n478_ = ~new_n472_ & new_n477_;
  assign new_n479_ = inp13 & new_n478_;
  assign otp17 = ~new_n463_ & ~new_n479_;
  assign new_n481_ = ~new_n214_ & new_n352_;
  assign new_n482_ = new_n214_ & ~new_n352_;
  assign new_n483_ = ~new_n481_ & ~new_n482_;
  assign new_n484_ = ~inp10 & ~new_n483_;
  assign new_n485_ = inp10 & new_n483_;
  assign new_n486_ = ~new_n484_ & ~new_n485_;
  assign new_n487_ = new_n68_ & new_n442_;
  assign new_n488_ = ~new_n486_ & new_n487_;
  assign new_n489_ = ~new_n325_ & ~new_n488_;
  assign new_n490_ = ~new_n68_ & new_n442_;
  assign new_n491_ = new_n486_ & new_n490_;
  assign new_n492_ = ~new_n327_ & ~new_n491_;
  assign otp16 = ~new_n489_ | ~new_n492_;
  assign new_n494_ = ~inp12 & inp9;
  assign new_n495_ = inp13 & new_n494_;
  assign new_n496_ = inp13 & ~inp11;
  assign new_n497_ = ~new_n217_ & new_n496_;
  assign new_n498_ = ~inp9 & ~new_n497_;
  assign new_n499_ = inp12 & ~new_n498_;
  assign new_n500_ = ~new_n138_ & ~new_n141_;
  assign new_n501_ = new_n138_ & new_n141_;
  assign new_n502_ = ~new_n500_ & ~new_n501_;
  assign new_n503_ = ~new_n499_ & ~new_n502_;
  assign new_n504_ = inp9 & ~new_n332_;
  assign new_n505_ = ~new_n503_ & ~new_n504_;
  assign new_n506_ = ~new_n495_ & ~new_n505_;
  assign new_n507_ = new_n217_ & new_n496_;
  assign new_n508_ = ~new_n334_ & ~new_n507_;
  assign new_n509_ = ~inp9 & ~new_n508_;
  assign new_n510_ = ~new_n144_ & ~new_n509_;
  assign new_n511_ = ~new_n506_ & ~new_n510_;
  assign otp15 = new_n331_ | new_n511_;
  assign new_n513_ = ~new_n81_ & ~new_n345_;
  assign new_n514_ = new_n71_ & new_n273_;
  assign new_n515_ = new_n144_ & ~new_n514_;
  assign new_n516_ = ~new_n513_ & new_n515_;
  assign new_n517_ = new_n81_ & ~new_n345_;
  assign new_n518_ = inp10 & new_n442_;
  assign new_n519_ = ~new_n144_ & ~new_n518_;
  assign new_n520_ = ~new_n517_ & new_n519_;
  assign new_n521_ = ~new_n516_ & ~new_n520_;
  assign otp14 = new_n343_ | new_n521_;
  assign new_n523_ = ~new_n279_ & new_n442_;
  assign new_n524_ = ~inp9 & ~new_n483_;
  assign new_n525_ = inp9 & new_n483_;
  assign new_n526_ = ~new_n524_ & ~new_n525_;
  assign new_n527_ = ~new_n353_ & ~new_n526_;
  assign new_n528_ = ~new_n68_ & ~new_n527_;
  assign new_n529_ = ~new_n523_ & new_n528_;
  assign new_n530_ = new_n279_ & new_n442_;
  assign new_n531_ = ~new_n353_ & new_n526_;
  assign new_n532_ = new_n68_ & ~new_n531_;
  assign new_n533_ = ~new_n530_ & new_n532_;
  assign new_n534_ = ~new_n529_ & ~new_n533_;
  assign otp13 = new_n362_ | new_n534_;
  assign new_n536_ = inp9 & inp6;
  assign new_n537_ = ~inp9 & ~inp6;
  assign new_n538_ = ~new_n536_ & ~new_n537_;
  assign new_n539_ = new_n173_ & new_n538_;
  assign new_n540_ = ~new_n173_ & ~new_n538_;
  assign new_n541_ = ~new_n539_ & ~new_n540_;
  assign new_n542_ = ~inp12 & ~new_n541_;
  assign new_n543_ = inp12 & new_n75_;
  assign new_n544_ = new_n141_ & ~new_n543_;
  assign new_n545_ = ~new_n542_ & new_n544_;
  assign new_n546_ = ~inp12 & new_n541_;
  assign new_n547_ = inp10 & new_n441_;
  assign new_n548_ = ~new_n141_ & ~new_n547_;
  assign new_n549_ = ~new_n546_ & new_n548_;
  assign new_n550_ = inp13 & ~new_n549_;
  assign new_n551_ = ~new_n545_ & new_n550_;
  assign otp12 = new_n373_ | new_n551_;
  assign new_n553_ = new_n279_ & new_n441_;
  assign new_n554_ = inp1 & new_n304_;
  assign new_n555_ = ~new_n553_ & ~new_n554_;
  assign new_n556_ = ~new_n71_ & ~new_n144_;
  assign new_n557_ = ~new_n352_ & ~new_n556_;
  assign new_n558_ = ~new_n71_ & new_n144_;
  assign new_n559_ = new_n352_ & ~new_n558_;
  assign new_n560_ = ~new_n557_ & ~new_n559_;
  assign new_n561_ = ~new_n84_ & ~new_n560_;
  assign new_n562_ = ~new_n352_ & ~new_n558_;
  assign new_n563_ = new_n352_ & ~new_n556_;
  assign new_n564_ = ~new_n562_ & ~new_n563_;
  assign new_n565_ = new_n84_ & ~new_n564_;
  assign new_n566_ = ~new_n561_ & ~new_n565_;
  assign new_n567_ = new_n437_ & new_n566_;
  assign new_n568_ = new_n555_ & ~new_n567_;
  assign new_n569_ = inp13 & ~new_n568_;
  assign new_n570_ = ~new_n84_ & ~new_n564_;
  assign new_n571_ = new_n84_ & ~new_n560_;
  assign new_n572_ = ~new_n570_ & ~new_n571_;
  assign new_n573_ = new_n495_ & new_n572_;
  assign new_n574_ = ~new_n375_ & ~new_n573_;
  assign otp11 = new_n569_ | ~new_n574_;
  assign new_n576_ = ~new_n402_ & ~new_n518_;
  assign otp10 = new_n400_ | ~new_n576_;
  assign new_n578_ = new_n285_ & new_n442_;
  assign otp9 = otp29 | new_n578_;
  assign otp8 = otp28 | new_n455_;
  assign new_n581_ = ~inp12 & inp7;
  assign new_n582_ = ~new_n65_ & ~new_n581_;
  assign new_n583_ = ~new_n459_ & new_n582_;
  assign new_n584_ = new_n458_ & ~new_n583_;
  assign new_n585_ = new_n441_ & ~new_n469_;
  assign new_n586_ = ~new_n494_ & ~new_n585_;
  assign new_n587_ = ~new_n141_ & ~new_n586_;
  assign new_n588_ = ~inp12 & new_n474_;
  assign new_n589_ = ~new_n476_ & ~new_n588_;
  assign new_n590_ = ~new_n587_ & new_n589_;
  assign new_n591_ = inp13 & ~new_n590_;
  assign otp7 = new_n584_ | new_n591_;
  assign new_n593_ = ~otp26 & ~new_n488_;
  assign otp6 = new_n491_ | ~new_n593_;
  assign new_n595_ = ~new_n334_ & ~new_n497_;
  assign new_n596_ = ~new_n138_ & new_n319_;
  assign new_n597_ = new_n138_ & new_n474_;
  assign new_n598_ = ~new_n596_ & ~new_n597_;
  assign new_n599_ = ~new_n595_ & ~new_n598_;
  assign new_n600_ = inp9 & new_n332_;
  assign new_n601_ = ~inp9 & new_n507_;
  assign new_n602_ = ~new_n600_ & ~new_n601_;
  assign new_n603_ = inp12 & ~new_n602_;
  assign new_n604_ = ~new_n495_ & ~new_n603_;
  assign new_n605_ = ~new_n144_ & ~new_n604_;
  assign new_n606_ = ~new_n599_ & ~new_n605_;
  assign otp5 = new_n331_ | ~new_n606_;
  assign new_n608_ = ~new_n513_ & new_n519_;
  assign new_n609_ = new_n515_ & ~new_n517_;
  assign new_n610_ = ~new_n608_ & ~new_n609_;
  assign otp4 = new_n343_ | new_n610_;
  assign new_n612_ = ~new_n68_ & ~new_n523_;
  assign new_n613_ = ~new_n531_ & new_n612_;
  assign new_n614_ = new_n68_ & ~new_n530_;
  assign new_n615_ = ~new_n527_ & new_n614_;
  assign new_n616_ = ~new_n613_ & ~new_n615_;
  assign otp3 = new_n362_ | new_n616_;
  assign new_n618_ = ~new_n542_ & new_n548_;
  assign new_n619_ = new_n544_ & ~new_n546_;
  assign new_n620_ = inp13 & ~new_n619_;
  assign new_n621_ = ~new_n618_ & new_n620_;
  assign otp2 = new_n373_ | new_n621_;
  assign new_n623_ = new_n437_ & new_n572_;
  assign new_n624_ = new_n555_ & ~new_n623_;
  assign new_n625_ = inp13 & ~new_n624_;
  assign new_n626_ = new_n495_ & new_n566_;
  assign new_n627_ = ~new_n375_ & ~new_n626_;
  assign otp1 = new_n625_ | ~new_n627_;
  assign otp0 = new_n429_ | ~new_n576_;
endmodule


